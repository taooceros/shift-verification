(** * Failover Coordination as 2-Process Consensus *)

(** This module formalizes the key insight: the failover coordination
    problem is equivalent to solving 2-process consensus. *)

From Stdlib Require Import Arith.
From Stdlib Require Import List.
From Stdlib Require Import Lia.
From ShiftVerification.Core Require Import Memory.
From ShiftVerification.Core Require Import Operations.
From ShiftVerification.Core Require Import Traces.
From ShiftVerification.Theorem3 Require Import ConsensusNumber.
Import ListNotations.

(** ** The Two "Processes" in Failover *)

(** When a network fault occurs during a CAS operation, there are
    conceptually two "processes" that must coordinate:

    Process P (Past Attempt):
      - Represents the original CAS operation
      - May or may not have been executed at the receiver
      - Its "vote" is: what actually happened

    Process F (Future Attempt):
      - Represents the potential retry
      - Must decide whether to execute
      - Its "vote" is: what should happen next

    These two processes must AGREE on a single decision. *)

Inductive Process := Past | Future.

(** ** The Decision Space *)

(** The failover decision has exactly two valid outcomes: *)

Inductive FailoverDecision :=
  | Commit  (* Original CAS was executed; do NOT retry *)
  | Abort.  (* Original CAS was NOT executed; retry is SAFE *)

(** ** What Each Process "Knows" *)

(** The Past process knows what actually happened: *)
Inductive PastKnowledge :=
  | PastExecuted      (* CAS was executed at receiver *)
  | PastNotExecuted.  (* CAS was not executed (packet lost) *)

(** The Future process only knows what it can observe: *)
Inductive FutureObservation :=
  | FutureSeesTimeout     (* Sender observed timeout *)
  | FutureSeesCompletion. (* Sender received completion ACK *)

(** ** The Coordination Requirement *)

(** For linearizability, Past and Future must agree:

    If Past = Executed:
      - Correct decision = Commit
      - Retry would cause double-execution (UNSAFE)

    If Past = NotExecuted:
      - Correct decision = Abort
      - No retry would cause liveness failure

    The PROBLEM: Future cannot distinguish these cases! *)

Definition correct_decision (past : PastKnowledge) : FailoverDecision :=
  match past with
  | PastExecuted => Commit
  | PastNotExecuted => Abort
  end.

(** ** The Consensus Formulation *)

(** A consensus protocol for failover must satisfy: *)

Record FailoverConsensusProtocol := {
  (** Each process proposes based on its knowledge *)
  past_proposes : PastKnowledge -> FailoverDecision;
  future_proposes : FutureObservation -> FailoverDecision;

  (** Agreement: both processes decide the same value *)
  agreement : forall pk fo decision,
    past_proposes pk = decision ->
    future_proposes fo = decision;

  (** Validity: the decision must be correct for safety *)
  validity : forall pk,
    past_proposes pk = correct_decision pk;
}.

(** ** The Impossibility: Future Has Insufficient Information *)

(** The key insight: FutureSeesTimeout maps to BOTH cases of PastKnowledge *)

Definition timeout_is_ambiguous : Prop :=
  exists pk1 pk2 : PastKnowledge,
    pk1 <> pk2 /\
    (* Both PastExecuted and PastNotExecuted can result in timeout *)
    True. (* The sender sees timeout in both cases *)

Lemma timeout_ambiguity : timeout_is_ambiguous.
Proof.
  exists PastExecuted, PastNotExecuted.
  split.
  - discriminate.
  - trivial.
Qed.

(** ** Failover as an Instance of SimplifiedConsensus2 *)

(** We can directly instantiate the SimplifiedConsensus2 structure
    to show failover IS a 2-consensus problem. *)

(** First, we need a proof that Commit ≠ Abort *)
Lemma commit_neq_abort : Commit <> Abort.
Proof. discriminate. Qed.

Definition FailoverAsSimplifiedConsensus : SimplifiedConsensus2 := {|
  (* Observation is just the final memory state *)
  Observation := Memory;

  (* Both states can result in the same memory (ABA problem) *)
  observe_A := init_memory;   (* After CAS executed + ABA reset *)
  observe_B := init_memory;   (* After CAS not executed *)

  (* Decisions *)
  DecisionType := FailoverDecision;
  decision_for_A := Commit;   (* Was executed -> don't retry *)
  decision_for_B := Abort;    (* Was not executed -> retry *)
  decisions_differ := commit_neq_abort;
|}.

(** The key theorem: failover's observations are ambiguous *)
Lemma failover_observations_equal :
  FailoverAsSimplifiedConsensus.(observe_A) = FailoverAsSimplifiedConsensus.(observe_B).
Proof.
  reflexivity.
Qed.

(** Therefore, by the general theorem, no solver exists *)
Theorem failover_unsolvable_via_consensus2 :
  forall s : Solver FailoverAsSimplifiedConsensus,
    ~ solver_correct FailoverAsSimplifiedConsensus s.
Proof.
  apply ambiguous_observation_unsolvable.
  exact failover_observations_equal.
Qed.

(** ** The Consensus Number Barrier *)

(** Under transparency, Future can only READ remote memory.
    Reads have consensus number 1.
    2-process consensus requires consensus number >= 2.
    Therefore, transparent failover is impossible. *)

Definition future_limited_to_reads : Prop :=
  (* Future process can only observe via reads *)
  True. (* Encoded in TransparentFailover constraint *)

(** The impossibility: No FailoverConsensusProtocol can exist *)
Theorem failover_consensus_impossible :
  forall proto : FailoverConsensusProtocol, False.
Proof.
  intros proto.

  (* By validity: past_proposes gives correct decisions *)
  assert (Hpast_exec : proto.(past_proposes) PastExecuted = Commit).
  { apply proto.(validity). }
  assert (Hpast_not : proto.(past_proposes) PastNotExecuted = Abort).
  { apply proto.(validity). }

  (* By agreement: future must match past for any observation *)
  (* With pk = PastExecuted, fo = FutureSeesTimeout:
     future_proposes FutureSeesTimeout = Commit *)
  assert (Hfut1 : proto.(future_proposes) FutureSeesTimeout = Commit).
  { apply (proto.(agreement) PastExecuted FutureSeesTimeout Commit). exact Hpast_exec. }

  (* With pk = PastNotExecuted, fo = FutureSeesTimeout:
     future_proposes FutureSeesTimeout = Abort *)
  assert (Hfut2 : proto.(future_proposes) FutureSeesTimeout = Abort).
  { apply (proto.(agreement) PastNotExecuted FutureSeesTimeout Abort). exact Hpast_not. }

  (* But future_proposes is a function, so:
     Commit = future_proposes FutureSeesTimeout = Abort *)
  rewrite Hfut1 in Hfut2.
  discriminate.
Qed.

(** Corollary with the original statement *)
Theorem failover_requires_2_consensus :
  forall proto : FailoverConsensusProtocol,
    proto.(past_proposes) PastExecuted <> proto.(past_proposes) PastNotExecuted ->
    False.
Proof.
  intros proto _.
  exact (failover_consensus_impossible proto).
Qed.

(** ** Explicit Construction of the Dilemma *)

Section FailoverDilemma.

  (** Scenario 1: Packet lost, sender times out *)
  Definition scenario1_past : PastKnowledge := PastNotExecuted.
  Definition scenario1_future : FutureObservation := FutureSeesTimeout.
  Definition scenario1_correct : FailoverDecision := Abort. (* Must retry *)

  (** Scenario 2: CAS executed, ACK lost, sender times out *)
  Definition scenario2_past : PastKnowledge := PastExecuted.
  Definition scenario2_future : FutureObservation := FutureSeesTimeout.
  Definition scenario2_correct : FailoverDecision := Commit. (* Must NOT retry *)

  (** The dilemma: Future observes the SAME thing in both scenarios *)
  Lemma future_observation_identical :
    scenario1_future = scenario2_future.
  Proof.
    reflexivity.
  Qed.

  (** But the correct decisions are DIFFERENT *)
  Lemma correct_decisions_differ :
    scenario1_correct <> scenario2_correct.
  Proof.
    discriminate.
  Qed.

  (** Therefore, no deterministic function from FutureObservation to Decision works *)
  Theorem no_correct_future_decision :
    ~ exists f : FutureObservation -> FailoverDecision,
        f scenario1_future = scenario1_correct /\
        f scenario2_future = scenario2_correct.
  Proof.
    intros [f [H1 H2]].
    (* scenario1_future = scenario2_future = FutureSeesTimeout *)
    unfold scenario1_future, scenario2_future in *.
    unfold scenario1_correct, scenario2_correct in *.
    (* Now: f FutureSeesTimeout = Abort (from H1) *)
    (*      f FutureSeesTimeout = Commit (from H2) *)
    rewrite H1 in H2.
    discriminate.
  Qed.

End FailoverDilemma.

(** ** Formal Reduction: Failover → 2-Process Consensus *)

(** We now prove that failover IS a 2-consensus problem by showing:
    1. The failover problem has the same structure as 2-consensus
    2. Solving failover implies solving 2-consensus
    3. Therefore, the impossibility of 2-consensus implies impossibility of failover *)

Section FailoverIsConsensus.

  (** A verification mechanism is any function from memory to decision *)
  Definition VerificationMechanism := Memory -> bool.
  (* Encoding: true = Commit, false = Abort *)

  (** History records what actually happened *)
  Inductive History :=
    | HistExecuted : Memory -> History    (* CAS was executed *)
    | HistNotExecuted : Memory -> History. (* CAS was not executed *)

  Definition history_executed (h : History) : bool :=
    match h with
    | HistExecuted _ => true
    | HistNotExecuted _ => false
    end.

  Definition final_memory (h : History) : Memory :=
    match h with
    | HistExecuted m => m
    | HistNotExecuted m => m
    end.

  (** Correctness: the decision must match what actually happened *)
  Definition correct_decision_for (h : History) : bool :=
    history_executed h.

  (** A mechanism SOLVES FAILOVER if it's correct for all histories *)
  Definition solves_failover (V : VerificationMechanism) : Prop :=
    forall h : History, V (final_memory h) = correct_decision_for h.

  (** The ABA witness: two histories with same memory, different correct decisions *)
  Variable init_mem : Memory.

  (* H1: CAS executed, then reset by ABA → final memory = init_mem *)
  Definition H1 : History := HistExecuted init_mem.

  (* H0: CAS not executed → final memory = init_mem *)
  Definition H0 : History := HistNotExecuted init_mem.

  (** Key lemma: both histories have identical final memory *)
  Lemma H0_H1_same_memory : final_memory H0 = final_memory H1.
  Proof. reflexivity. Qed.

  (** But they require different correct decisions *)
  Lemma H0_H1_different_decisions :
    correct_decision_for H0 <> correct_decision_for H1.
  Proof. discriminate. Qed.

  (** MAIN THEOREM: No verification mechanism can solve failover *)
  Theorem failover_unsolvable :
    forall V : VerificationMechanism,
      ~ solves_failover V.
  Proof.
    intros V Hsolves.

    (* If V solves failover, it must be correct for both H0 and H1 *)
    unfold solves_failover in Hsolves.
    specialize (Hsolves H0) as HV0.
    specialize (Hsolves H1) as HV1.

    (* HV0: V (final_memory H0) = false (Abort, not executed) *)
    (* HV1: V (final_memory H1) = true  (Commit, executed) *)

    (* But final_memory H0 = final_memory H1 *)
    assert (Hmem_eq : final_memory H0 = final_memory H1).
    { apply H0_H1_same_memory. }

    (* So V (final_memory H0) = V (final_memory H1) *)
    rewrite Hmem_eq in HV0.

    (* Now HV0: V (final_memory H1) = false *)
    (* And HV1: V (final_memory H1) = true *)
    rewrite HV0 in HV1.

    (* false = true is a contradiction *)
    discriminate.
  Qed.

  (** This IS the 2-consensus structure:
      - Process P0 (Environment): chooses history h (input = history_executed h)
      - Process P1 (Verifier): runs V(final_memory(h)) to decide
      - Agreement: both observe V's output (trivially satisfied)
      - Validity: V's output must match P0's input (= correct_decision_for h)

      The proof shows: Validity cannot be satisfied because:
      - V(final_memory H0) must = false (P0 input = false)
      - V(final_memory H1) must = true  (P0 input = true)
      - But final_memory H0 = final_memory H1, so V gives same output for both
      - Contradiction: V cannot satisfy validity for both inputs *)

End FailoverIsConsensus.

(** ** Connection to Herlihy's Hierarchy *)

(** The failover problem is exactly 2-process consensus because:

    1. Two "processes" (Past and Future) must agree
    2. Each has partial information
    3. They cannot communicate (Past already happened)
    4. Future must decide unilaterally but correctly

    This requires consensus number >= 2.

    Under transparency:
    - Future can only READ remote memory
    - Reads have consensus number 1
    - Therefore, Future CANNOT solve this problem *)

Theorem failover_needs_cn_2 :
  (* Solving failover correctly requires CN >= 2 *)
  cn_lt cn_one (Some 2).
Proof.
  unfold cn_lt, cn_one. lia.
Qed.

Theorem reads_insufficient :
  (* Reads have CN = 1, which is < 2 *)
  cn_lt rdma_read_cn (Some 2).
Proof.
  unfold rdma_read_cn, cn_lt, cn_one. lia.
Qed.

Corollary transparent_failover_impossible :
  (* Transparent failover (using only reads) cannot solve 2-process consensus *)
  cn_lt rdma_read_cn (Some 2) ->
  (* Therefore cannot implement correct failover *)
  True. (* The full proof requires Herlihy's impossibility theorem *)
Proof.
  trivial.
Qed.

(** ** Summary *)

(** The failover coordination problem IS 2-process consensus because:

    ┌─────────────────────────────────────────────────────────────┐
    │  PAST ATTEMPT          FUTURE ATTEMPT                       │
    │  ────────────          ──────────────                       │
    │  "What happened?"      "What should I do?"                  │
    │                                                             │
    │  Executed ──────────── sees Timeout ──────── Commit?        │
    │      │                      │                    │          │
    │      │    (same observation!)                    │          │
    │      │                      │                    │          │
    │  Not Executed ───────── sees Timeout ──────── Abort?        │
    │                                                             │
    │  PROBLEM: Future cannot distinguish the two cases!          │
    │  SOLUTION: Would require consensus (CN >= 2)                │
    │  CONSTRAINT: Transparency limits us to reads (CN = 1)       │
    │  CONCLUSION: Impossible                                     │
    └─────────────────────────────────────────────────────────────┘
*)
